class top_sqr extends uvm_sequencer;
write_sqr write_sqr_i;
read_sqr read_sqr_i;
`uvm_component_utils(top_sqr)
`NEW_COMP

endclass
